/*
This module was out generated using maasm, MiniAlu's assembler
report any bug to javinachop@gmail.com

maasm is distributed under GNU GPL see <http://www.gnu.org/licenses/>
*/
`ifndef ROM_A
`define ROM_A


`timescale 1ns / 1ps
module ROM(
	   input wire [31:0] iAddress,
	   output reg [31:0] oInstruction
	   );
 always @ ( iAddress )
     begin
	case (iAddress)
          
           0: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           1: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           2: oInstruction = 32'b00001011101000000000000000000000; // addiu $sp $0 0
          
           3: oInstruction = 32'b00111111101111011000000000000000; // sll $sp $sp 16
          
           4: oInstruction = 32'b00110111101000000000000100111100; // ori $sp $0 316
          
           5: oInstruction = 32'b00001011110000000000000000000000; // addiu $fp $0 0
          
           6: oInstruction = 32'b00111111110111101000000000000000; // sll $fp $fp 16
          
           7: oInstruction = 32'b00110111110000000000000100111100; // ori $fp $0 316
          
           8: oInstruction = 32'b01011100000000000000000010011111; // j main
          
           9: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           10: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           11: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           12: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           13: oInstruction = 32'b00010111101111010000000000101000; // subi $sp $sp -40
          
           14: oInstruction = 32'b10010011111111010000000000100100; // sw $31 36 $sp
          
           15: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           16: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           17: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           18: oInstruction = 32'b10010011110111010000000000100000; // sw $fp 32 $sp
          
           19: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           20: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           21: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           22: oInstruction = 32'b00001111110111010000000000000000; // move $fp $sp
          
           23: oInstruction = 32'b10010000100111100000000000101000; // sw $4 40 $fp
          
           24: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           25: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           26: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           27: oInstruction = 32'b10010000101111100000000000101100; // sw $5 44 $fp
          
           28: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           29: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           30: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           31: oInstruction = 32'b10001100011111100000000000101100; // lw $3 44 $fp
          
           32: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           33: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           34: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           35: oInstruction = 32'b00001000010000000000000000000000; // addiu $2 $0 0
          
           36: oInstruction = 32'b00111100010000101000000000000000; // sll $2 $2 16
          
           37: oInstruction = 32'b00110100010000000000000000000001; // ori $2 $0 1
          
           38: oInstruction = 32'b10000000011000100000000001001010; // bne $3 $2 $L2
          
           39: oInstruction = 32'b00001000010000000000000000000000; // addiu $2 $0 0
          
           40: oInstruction = 32'b00111100010000101000000000000000; // sll $2 $2 16
          
           41: oInstruction = 32'b00110100010000000000000000000001; // ori $2 $0 1
          
           42: oInstruction = 32'b10010000010111100000000000010100; // sw $2 20 $fp
          
           43: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           44: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           45: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           46: oInstruction = 32'b00001000010000000000000000000000; // addiu $2 $0 0
          
           47: oInstruction = 32'b00111100010000101000000000000000; // sll $2 $2 16
          
           48: oInstruction = 32'b00110100010000000000000000000010; // ori $2 $0 2
          
           49: oInstruction = 32'b10010000010111100000000000011000; // sw $2 24 $fp
          
           50: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           51: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           52: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           53: oInstruction = 32'b10001100010111100000000000101000; // lw $2 40 $fp
          
           54: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           55: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           56: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           57: oInstruction = 32'b10001100100111100000000000010100; // lw $4 20 $fp
          
           58: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           59: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           60: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           61: oInstruction = 32'b10001100011111100000000000011000; // lw $3 24 $fp
          
           62: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           63: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           64: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           65: oInstruction = 32'b10010000100000100000000000000000; // sw $4 0 $2
          
           66: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           67: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           68: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           69: oInstruction = 32'b10010000011000100000000000000100; // sw $3 4 $2
          
           70: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           71: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           72: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           73: oInstruction = 32'b01011100000000000000000010010000; // b $L1
          
           74: oInstruction = 32'b10001100010111100000000000101100; // lw $2 44 $fp
          
           75: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           76: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           77: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           78: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           79: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           80: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           81: oInstruction = 32'b00010100011000100000000000000001; // subi $3 $2 -1
          
           82: oInstruction = 32'b00001000010111100000000000010100; // addiu $2 $fp 20
          
           83: oInstruction = 32'b00001100101000110000000000000000; // move $5 $3
          
           84: oInstruction = 32'b00001100100000100000000000000000; // move $4 $2
          
           85: oInstruction = 32'b01111000000000000000000000001101; // jal fibonacci
          
           86: oInstruction = 32'b10001100010111100000000000011000; // lw $2 24 $fp
          
           87: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           88: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           89: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           90: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           91: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           92: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           93: oInstruction = 32'b10010000010111100000000000010000; // sw $2 16 $fp
          
           94: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           95: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           96: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           97: oInstruction = 32'b10001100011111100000000000011000; // lw $3 24 $fp
          
           98: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           99: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           100: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           101: oInstruction = 32'b10001100010111100000000000010100; // lw $2 20 $fp
          
           102: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           103: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           104: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           105: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           106: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           107: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           108: oInstruction = 32'b00001100010000110001000000000000; // addu $2 $3 $2
          
           109: oInstruction = 32'b10010000010111100000000000011000; // sw $2 24 $fp
          
           110: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           111: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           112: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           113: oInstruction = 32'b10001100010111100000000000010000; // lw $2 16 $fp
          
           114: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           115: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           116: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           117: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           118: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           119: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           120: oInstruction = 32'b10010000010111100000000000010100; // sw $2 20 $fp
          
           121: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           122: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           123: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           124: oInstruction = 32'b10001100010111100000000000101000; // lw $2 40 $fp
          
           125: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           126: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           127: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           128: oInstruction = 32'b10001100100111100000000000010100; // lw $4 20 $fp
          
           129: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           130: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           131: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           132: oInstruction = 32'b10001100011111100000000000011000; // lw $3 24 $fp
          
           133: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           134: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           135: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           136: oInstruction = 32'b10010000100000100000000000000000; // sw $4 0 $2
          
           137: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           138: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           139: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           140: oInstruction = 32'b10010000011000100000000000000100; // sw $3 4 $2
          
           141: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           142: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           143: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           144: oInstruction = 32'b10001100010111100000000000101000; // lw $2 40 $fp
          
           145: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           146: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           147: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           148: oInstruction = 32'b00001111101111100000000000000000; // move $sp $fp
          
           149: oInstruction = 32'b10001111111111010000000000100100; // lw $31 36 $sp
          
           150: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           151: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           152: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           153: oInstruction = 32'b10001111110111010000000000100000; // lw $fp 32 $sp
          
           154: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           155: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           156: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           157: oInstruction = 32'b00001011101111010000000000101000; // addiu $sp $sp 40
          
           158: oInstruction = 32'b01100000000000001111100000000000; // jr $ra
          
           159: oInstruction = 32'b00010111101111010000000000101000; // subi $sp $sp -40
          
           160: oInstruction = 32'b10010011111111010000000000100100; // sw $31 36 $sp
          
           161: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           162: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           163: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           164: oInstruction = 32'b10010011110111010000000000100000; // sw $fp 32 $sp
          
           165: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           166: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           167: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           168: oInstruction = 32'b00001111110111010000000000000000; // move $fp $sp
          
           169: oInstruction = 32'b00001000010000000000000000000000; // addiu $2 $0 0
          
           170: oInstruction = 32'b00111100010000101000000000000000; // sll $2 $2 16
          
           171: oInstruction = 32'b00110100010000000000000000000010; // ori $2 $0 2
          
           172: oInstruction = 32'b10010000010111100000000000010000; // sw $2 16 $fp
          
           173: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           174: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           175: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           176: oInstruction = 32'b01011100000000000000000011001100; // b $L6
          
           177: oInstruction = 32'b00001000010111100000000000010100; // addiu $2 $fp 20
          
           178: oInstruction = 32'b10001100101111100000000000010000; // lw $5 16 $fp
          
           179: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           180: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           181: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           182: oInstruction = 32'b00001100100000100000000000000000; // move $4 $2
          
           183: oInstruction = 32'b01111000000000000000000000001101; // jal fibonacci
          
           184: oInstruction = 32'b10001100010111100000000000011000; // lw $2 24 $fp
          
           185: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           186: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           187: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           188: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           189: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           190: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           191: oInstruction = 32'b10010100000000100000000000000000; // led $2
          
           192: oInstruction = 32'b10001100010111100000000000010000; // lw $2 16 $fp
          
           193: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           194: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           195: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           196: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           197: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           198: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           199: oInstruction = 32'b00001000010000100000000000000001; // addiu $2 $2 1
          
           200: oInstruction = 32'b10010000010111100000000000010000; // sw $2 16 $fp
          
           201: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           202: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           203: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           204: oInstruction = 32'b10001100010111100000000000010000; // lw $2 16 $fp
          
           205: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           206: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           207: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           208: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           209: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           210: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           211: oInstruction = 32'b00101100010000100000000000000110; // slti $2 $2 6
          
           212: oInstruction = 32'b10000000010000000000000010110001; // bne $2 $0 $L7
          
           213: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           214: oInstruction = 32'b00001111101111100000000000000000; // move $sp $fp
          
           215: oInstruction = 32'b10001111111111010000000000100100; // lw $31 36 $sp
          
           216: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           217: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           218: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           219: oInstruction = 32'b10001111110111010000000000100000; // lw $fp 32 $sp
          
           220: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           221: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           222: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           223: oInstruction = 32'b00001011101111010000000000101000; // addiu $sp $sp 40
          
           224: oInstruction = 32'b01011100000000000000000010011111; // j main
          
           225: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           226: oInstruction = 32'b00000000000000000000000000000000; // nop
          
           227: oInstruction = 32'b00000000000000000000000000000000; // nop
          
	  default:
	    oInstruction = { 4'b0010 ,  24'b10101010 };		//NOP
	endcase
     end

endmodule
`endif //ROM_A